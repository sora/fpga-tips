module testbench;
	initial begin
		$display("Hello World");
		$display("Hello World");
		$display("Hello World");
		$display("Hello World");

		$finish;
	end
endmodule
